module PC_Adder(
    IM_busy,
    DM_busy,
    Flush,
    JALR,
    U_AUIPC,
    PC,
    imm32,
    Data_rs1,
    New_PC,
    PC_branch,
    PCAdd4
);

input   IM_busy, DM_busy, Flush, JALR, U_AUIPC;
input   [31:0]  PC, imm32, Data_rs1;    
output  [31:0]  New_PC, PC_branch, PCAdd4;

wire    [31:0]  choice, PC_branch, PCAdd4;

assign  choice = (~JALR | U_AUIPC)? (PC - 32'd4) : Data_rs1;
assign  PC_branch = choice + imm32 ;
assign  PCAdd4 = PC+32'd4;
//assign  New_PC = (IM_busy)? PC : ((Flush)? PC_branch : PCAdd4);
//assign  New_PC = (IM_busy | DM_busy)? PC : ((Flush)? PC_branch : PCAdd4);
assign  New_PC = (Flush)? PC_branch : ((IM_busy | DM_busy)? PC : PCAdd4);

endmodule
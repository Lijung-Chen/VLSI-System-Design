//stalling pipeline
module  Hazard_detection(
    Branch,
    ID_EX_MemRead,
    ID_EX_Rd,
    EX_MEM_MemRead,
    EX_MEM_Rd,
    ID_EX_RegWrite,
    IF_ID_RS1,
    IF_ID_RS2,
    ID_EX_MULtype,
    mul_finish,
    IF_ID_Write,
    PC_Write,
    Stall
);

input       Branch, ID_EX_MemRead, EX_MEM_MemRead, ID_EX_RegWrite, mul_finish;
input       [1:0]ID_EX_MULtype;
input       [4:0]ID_EX_Rd, EX_MEM_Rd, IF_ID_RS1, IF_ID_RS2;
output  reg IF_ID_Write, PC_Write, Stall;

always@(*)begin
    if(ID_EX_MemRead && (ID_EX_Rd == IF_ID_RS1 || ID_EX_Rd == IF_ID_RS2)) begin //lw+R
        IF_ID_Write = 1'b0;
        PC_Write = 1'b0;
        Stall = 1'b1;
    end
    else if(Branch && EX_MEM_MemRead && (EX_MEM_Rd == IF_ID_RS1 || EX_MEM_Rd == IF_ID_RS2)) begin   //lw+B
        IF_ID_Write = 1'b0;
        PC_Write = 1'b0;
        Stall = 1'b1;
    end
    else if(Branch && ID_EX_RegWrite && (ID_EX_Rd == IF_ID_RS1 || ID_EX_Rd == IF_ID_RS2)) begin   //R+B
        IF_ID_Write = 1'b0;
        PC_Write = 1'b0;
        Stall = 1'b1;
    end
    else if(ID_EX_MULtype != 2'd0 && !mul_finish) begin
        IF_ID_Write = 1'b0;
        PC_Write = 1'b0;
        Stall = 1'b1;
    end
    else begin
        IF_ID_Write = 1'b1;
        PC_Write = 1'b1;
        Stall = 1'b0;
    end
end

endmodule